module e2q3(a,b,c,rw,rd,alu,mr,mw,mtor,br,j);
input a,b,c;
output rw,rd,alu,mr,mw,mtor,br,j;


endmodule 
