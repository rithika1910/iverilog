module mux4x1_using_2x1mux_tb();
reg s0,s1,i0,i1,i2,i3;
wire y;

mux4x1_using_2x1mux muxtb4x1(i0, i1, i2, i3, s0, s1, y);
initial
begin
  $display(" | S0 | S1 | I0 | I1 | I2 | I3 | Y | ");
  $monitor(" | %b  | %b  | %b  | %b  | %b  | %b  | %b | ",s0,s1,i0,i1,i2,i3,y);
  s0 = 0; s1 = 0; i0 = 0; i1 = 0; i2 = 0; i3 = 0 ; #10;
  s0 = 0; s1 = 0; i0 = 0; i1 = 0; i2 = 0; i3 = 1 ; #10;
  s0 = 0; s1 = 0; i0 = 0; i1 = 0; i2 = 1; i3 = 0 ; #10;
  s0 = 0; s1 = 0; i0 = 0; i1 = 0; i2 = 1; i3 = 1 ; #10;
  s0 = 0; s1 = 0; i0 = 0; i1 = 1; i2 = 0; i3 = 0 ; #10;
  s0 = 0; s1 = 0; i0 = 0; i1 = 1; i2 = 0; i3 = 1 ; #10;
  s0 = 0; s1 = 0; i0 = 0; i1 = 1; i2 = 1; i3 = 0 ; #10;
  s0 = 0; s1 = 0; i0 = 0; i1 = 1; i2 = 1; i3 = 1 ; #10;
  s0 = 0; s1 = 0; i0 = 1; i1 = 0; i2 = 0; i3 = 0 ; #10;
  s0 = 0; s1 = 0; i0 = 1; i1 = 0; i2 = 0; i3 = 1 ; #10;
  s0 = 0; s1 = 0; i0 = 1; i1 = 0; i2 = 1; i3 = 0 ; #10;
  s0 = 0; s1 = 0; i0 = 1; i1 = 0; i2 = 1; i3 = 1 ; #10;
  s0 = 0; s1 = 0; i0 = 1; i1 = 1; i2 = 0; i3 = 0 ; #10;
  s0 = 0; s1 = 0; i0 = 1; i1 = 1; i2 = 0; i3 = 1 ; #10;
  s0 = 0; s1 = 0; i0 = 1; i1 = 1; i2 = 1; i3 = 0 ; #10;
  s0 = 0; s1 = 0; i0 = 1; i1 = 1; i2 = 1; i3 = 1 ; #10;

  s0 = 0; s1 = 1; i0 = 0; i1 = 0; i2 = 0; i3 = 0 ; #10;
  s0 = 0; s1 = 1; i0 = 0; i1 = 0; i2 = 0; i3 = 1 ; #10;
  s0 = 0; s1 = 1; i0 = 0; i1 = 0; i2 = 1; i3 = 0 ; #10;
  s0 = 0; s1 = 1; i0 = 0; i1 = 0; i2 = 1; i3 = 1 ; #10;
  s0 = 0; s1 = 1; i0 = 0; i1 = 1; i2 = 0; i3 = 0 ; #10;
  s0 = 0; s1 = 1; i0 = 0; i1 = 1; i2 = 0; i3 = 1 ; #10;
  s0 = 0; s1 = 1; i0 = 0; i1 = 1; i2 = 1; i3 = 0 ; #10;
  s0 = 0; s1 = 1; i0 = 0; i1 = 1; i2 = 1; i3 = 1 ; #10;
  s0 = 0; s1 = 1; i0 = 1; i1 = 0; i2 = 0; i3 = 0 ; #10;
  s0 = 0; s1 = 1; i0 = 1; i1 = 0; i2 = 0; i3 = 1 ; #10;
  s0 = 0; s1 = 1; i0 = 1; i1 = 0; i2 = 1; i3 = 0 ; #10;
  s0 = 0; s1 = 1; i0 = 1; i1 = 0; i2 = 1; i3 = 1 ; #10;
  s0 = 0; s1 = 1; i0 = 1; i1 = 1; i2 = 0; i3 = 0 ; #10;
  s0 = 0; s1 = 1; i0 = 1; i1 = 1; i2 = 0; i3 = 1 ; #10;
  s0 = 0; s1 = 1; i0 = 1; i1 = 1; i2 = 1; i3 = 0 ; #10;
  s0 = 0; s1 = 1; i0 = 1; i1 = 1; i2 = 1; i3 = 1 ; #10;

  s0 = 1; s1 = 0; i0 = 0; i1 = 0; i2 = 0; i3 = 0 ; #10;
  s0 = 1; s1 = 0; i0 = 0; i1 = 0; i2 = 0; i3 = 1 ; #10;
  s0 = 1; s1 = 0; i0 = 0; i1 = 0; i2 = 1; i3 = 0 ; #10;
  s0 = 1; s1 = 0; i0 = 0; i1 = 0; i2 = 1; i3 = 1 ; #10;
  s0 = 1; s1 = 0; i0 = 0; i1 = 1; i2 = 0; i3 = 0 ; #10;
  s0 = 1; s1 = 0; i0 = 0; i1 = 1; i2 = 0; i3 = 1 ; #10;
  s0 = 1; s1 = 0; i0 = 0; i1 = 1; i2 = 1; i3 = 0 ; #10;
  s0 = 1; s1 = 0; i0 = 0; i1 = 1; i2 = 1; i3 = 1 ; #10;
  s0 = 1; s1 = 0; i0 = 1; i1 = 0; i2 = 0; i3 = 0 ; #10;
  s0 = 1; s1 = 0; i0 = 1; i1 = 0; i2 = 0; i3 = 1 ; #10;
  s0 = 1; s1 = 0; i0 = 1; i1 = 0; i2 = 1; i3 = 0 ; #10;
  s0 = 1; s1 = 0; i0 = 1; i1 = 0; i2 = 1; i3 = 1 ; #10;
  s0 = 1; s1 = 0; i0 = 1; i1 = 1; i2 = 0; i3 = 0 ; #10;
  s0 = 1; s1 = 0; i0 = 1; i1 = 1; i2 = 0; i3 = 1 ; #10;
  s0 = 1; s1 = 0; i0 = 1; i1 = 1; i2 = 1; i3 = 0 ; #10;
  s0 = 1; s1 = 0; i0 = 1; i1 = 1; i2 = 1; i3 = 1 ; #10;

  s0 = 1; s1 = 1; i0 = 0; i1 = 0; i2 = 0; i3 = 0 ; #10;
  s0 = 1; s1 = 1; i0 = 0; i1 = 0; i2 = 0; i3 = 1 ; #10;
  s0 = 1; s1 = 1; i0 = 0; i1 = 0; i2 = 1; i3 = 0 ; #10;
  s0 = 1; s1 = 1; i0 = 0; i1 = 0; i2 = 1; i3 = 1 ; #10;
  s0 = 1; s1 = 1; i0 = 0; i1 = 1; i2 = 0; i3 = 0 ; #10;
  s0 = 1; s1 = 1; i0 = 0; i1 = 1; i2 = 0; i3 = 1 ; #10;
  s0 = 1; s1 = 1; i0 = 0; i1 = 1; i2 = 1; i3 = 0 ; #10;
  s0 = 1; s1 = 1; i0 = 0; i1 = 1; i2 = 1; i3 = 1 ; #10;
  s0 = 1; s1 = 1; i0 = 1; i1 = 0; i2 = 0; i3 = 0 ; #10;
  s0 = 1; s1 = 1; i0 = 1; i1 = 0; i2 = 0; i3 = 1 ; #10;
  s0 = 1; s1 = 1; i0 = 1; i1 = 0; i2 = 1; i3 = 0 ; #10;
  s0 = 1; s1 = 1; i0 = 1; i1 = 0; i2 = 1; i3 = 1 ; #10;
  s0 = 1; s1 = 1; i0 = 1; i1 = 1; i2 = 0; i3 = 0 ; #10;
  s0 = 1; s1 = 1; i0 = 1; i1 = 1; i2 = 0; i3 = 1 ; #10;
  s0 = 1; s1 = 1; i0 = 1; i1 = 1; i2 = 1; i3 = 0 ; #10;
  s0 = 1; s1 = 1; i0 = 1; i1 = 1; i2 = 1; i3 = 1 ; #10;
  $finish;
end
endmodule
